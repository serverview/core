<!DOCTYPE html>
<html lang="en">
<head>
    <meta charset="UTF-8">
    <meta name="viewport" content="width=device-width, initial-scale=1.0">
    <title>Hello from SVH</title>
</head>
<body>
    <p>Hi from SVH on version <system get="version"></system>.</p>
</body>
</html>